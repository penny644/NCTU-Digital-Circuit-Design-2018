module Lab2_BCD_7segment_decoder_behavior (A,D);
	output reg [6:0] A;
	input [3:0] D;
	always@(*)
	 begin 
	  A[0]=!D[3]&(D[1])|(!D[3])&D[2]&D[0]|D[3]&(!D[2])&!D[1]|(!D[2])&(!D[1])&(!D[0]);
	  A[1]=(!D[3])&(!D[2])|D[3]&(!D[2])&(!D[1])|(!D[3])&(!D[1])&(!D[0])|(!D[3])&D[1]&D[0];
	  A[2]=(!D[2])&(!D[1])|(!D[3])&D[2]|(!D[3])&D[0];
	  A[3]=(!D[3])&D[2]&(!D[1])&D[0]|D[3]&(!D[2])&(!D[1])|(!D[2])&(!D[1])&(!D[0])|(!D[3])&(!D[2])&D[1]|(!D[3])&D[1]&(!D[0]);
	  A[4]=(!D[3])&D[1]&(!D[0])|(!D[2])&(!D[1])&(!D[0]);
	  A[5]=D[3]&(!D[2])&(!D[1])|(!D[3])&D[2]&(!D[1])|(!D[3])&D[2]&(!D[0])|(!D[3])&(!D[1])&(!D[0]);
	  A[6]=D[3]&(!D[2])&(!D[1])|(!D[3])&D[2]&(!D[1])|(!D[3])&(!D[2])&D[1]|(!D[3])&D[1]&(!D[0]);
	 end
endmodule 
